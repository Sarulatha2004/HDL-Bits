module top_module ( input [1:0] A, input [1:0] B, output z ); 
    assign f = ~x3&x2 | x3&x1;

endmodule
